/*
 *  Write on positive clock edge
 *  Asynchronous read
 *
 *  Currently supports maximum of 64 instructions
 */

module instr_mem (
    input logic clk,
    input logic [9:0] read_addr,
    input logic [9:0] write_addr,
    input logic [31:0] write_instr,
    input logic write_en,

    output logic [31:0] read_instr
);

// Hard coded part of instruction memory containing
// the following common programs:
// 1. Reset frame buffer (fill with white)
// 2. Display horizontal white bars (used for top and bottom)
// 3. Display frame buffer
const logic [31:0] fixed_instrs [0:411] = {
    // Program 1: reset frame buffer
    // Starting address: 0d512
    32'h2001a824,
    32'h00018084,
    32'h80000480,
    32'h20040084,
    32'h80000480,
    32'h20040084,
    32'h80000480,
    32'h20040084,
    32'h80000480,
    32'h20040084,
    32'h80000480,
    32'h20040084,
    32'h80000480,
    32'h20040084,
    32'h80000480,
    32'h20040084,
    32'h80000480,
    32'h20040084,
    32'h80000480,
    32'h20040084,
    32'h80000480,
    32'h20040084,
    32'h80000480,
    32'h20040084,
    32'h80000480,
    32'h20040084,
    32'h80000480,
    32'h20040084,
    32'h80000480,
    32'h20040084,
    32'h80000480,
    32'h20040084,
    32'h80000480,
    32'h20040084,
    32'h80000480,
    32'h20040084,
    32'h80000480,
    32'h20040084,
    32'h80000480,
    32'h20040084,
    32'h80000480,
    32'h20040084,
    32'h80000480,
    32'h20040084,
    32'h80000480,
    32'h20040084,
    32'h80000480,
    32'h20040084,
    32'h80000480,
    32'h20040084,
    32'h80000480,
    32'h20040084,
    32'h80000480,
    32'h20040084,
    32'h80000480,
    32'h20040084,
    32'h80000480,
    32'h20040084,
    32'h80000480,
    32'h20040084,
    32'h80000480,
    32'h20040084,
    32'h80000480,
    32'h20040084,
    32'h80000480,
    32'h20040084,
    32'h80000480,
    32'h20040084,
    32'h80000480,
    32'h20040084,
    32'h80000480,
    32'h20040084,
    32'h80000480,
    32'h20040084,
    32'h80000480,
    32'h20040084,
    32'h80000480,
    32'h20040084,
    32'h80000480,
    32'h20040084,
    32'h80000480,
    32'h20040084,
    32'h80000480,
    32'h20040084,
    32'h80000480,
    32'h20040084,
    32'h80000480,
    32'h20040084,
    32'h80000480,
    32'h20040084,
    32'h80000480,
    32'h20040084,
    32'h80000480,
    32'h20040084,
    32'h80000480,
    32'h20040084,
    32'h80000480,
    32'h20040084,
    32'h80000480,
    32'h20040084,
    32'h80000480,
    32'h20040084,
    32'h80000480,
    32'h20040084,
    32'h80000480,
    32'h20040084,
    32'h80000480,
    32'h20040084,
    32'h80000480,
    32'h20040084,
    32'h80000480,
    32'h20040084,
    32'h80000480,
    32'h20040084,
    32'h80000480,
    32'h20040084,
    32'h80000480,
    32'h20040084,
    32'h80000480,
    32'h20040084,
    32'h80000480,
    32'h20040084,
    32'h80000480,
    32'h20040084,
    32'h80000480,
    32'h20040084,
    32'h80000480,
    32'h20040084,
    32'h80000480,
    32'h20040084,
    32'he0001c00,

    // Program 2: display horizontal white bar
    // Starting address: 0d643
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'he0001c00,

    // Program 3: display frame buffer
    // Starting address: 0d852
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'h20079c25,
    32'h2001a8a5,
    32'h000180a5,
    32'h20022c24,
    32'h2004a884,
    32'h00028084,
    32'h80000086,
    32'h20010007,
    32'h30000007,
    32'h000074c0,
    32'h20008488,
    32'h90000106,
    32'h100074c0,
    32'h21000488,
    32'h90000106,
    32'h100074c0,
    32'h21008488,
    32'h90000106,
    32'h2000f0e0,
    32'hc00000c0,
    32'h20400084,
    32'h80000086,
    32'h20010008,
    32'h30000008,
    32'h000074c0,
    32'h20008487,
    32'h900000e6,
    32'h100074c0,
    32'h21000487,
    32'h900000e6,
    32'h100074c0,
    32'h21008487,
    32'h900000e6,
    32'h2000f100,
    32'hc00000c0,
    32'h20400084,
    32'h80000086,
    32'h20010007,
    32'h30000007,
    32'h000074c0,
    32'h20008488,
    32'h90000106,
    32'h100074c0,
    32'h21000488,
    32'h90000106,
    32'h100074c0,
    32'h21008488,
    32'h90000106,
    32'h2000f0e0,
    32'hc00000c0,
    32'h20400084,
    32'h80000086,
    32'h20010008,
    32'h30000008,
    32'h000074c0,
    32'h20008487,
    32'h900000e6,
    32'h100074c0,
    32'h21000487,
    32'h900000e6,
    32'h100074c0,
    32'h21008487,
    32'h900000e6,
    32'h2000f100,
    32'hc00000c0,
    32'hc0000000,
    32'hc0000000,
    32'hc0000000,
    32'he0001c00
};

// 256-word programmable instruction memory
// Starts at address 0d0
logic [31:0] programmable_instrs [0:511];

always_comb begin
    read_instr = read_addr < 10'd512 ? programmable_instrs[read_addr[8:0]]
                                     : fixed_instrs[read_addr[8:0]];
end

always_ff @(posedge clk) begin
    if (write_en && write_addr < 10'd512) begin
        programmable_instrs[write_addr[8:0]] <= write_instr;
    end
end

endmodule
